library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constantesProcessador.all;

entity memoriaROM is

   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataROMWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataROMWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
        -- Inicializa os endereços: 
		   tmp(0) := "1001100000000000";
			tmp(1) := "1001100100000000";
			tmp(2) := "1001101000000000";
			tmp(3) := "1001101100000000";
			tmp(4) := "1001110000000000";
			tmp(5) := "1001110100000000";
			tmp(6) := "1001111000000000";
			tmp(7) := "1001111100000000";
			tmp(8) := "0000110000000000";
			tmp(9) := "0000000001000010";
			tmp(10) := "0000000101000011";
			tmp(11) := "1010000000000001";
			tmp(12) := "0001100000010000";
			tmp(13) := "1010000100000001";
			tmp(14) := "0001100000100010";
			tmp(15) := "0001000000001001";
			tmp(16) := "0000001001000001";
			tmp(17) := "1010001000000001";
			tmp(18) := "0001100000011000";
			tmp(19) := "1010001000000010";
			tmp(20) := "0001100000011111";
			tmp(21) := "1010001000000011";
			tmp(22) := "0001100000011010";
			tmp(23) := "0001000000011100";
			tmp(24) := "0000001101000000";
			tmp(25) := "0001000000001001";
			tmp(26) := "0000010001000000";
			tmp(27) := "0001000000001001";
			tmp(28) := "0000010101000000";
			tmp(29) := "0000100000001101";
			tmp(30) := "0001000000001001";
			tmp(31) := "0000011001000000";
			tmp(32) := "0000100000010110";
			tmp(33) := "0001000000001001";
			tmp(34) := "0000001001000000";
			tmp(35) := "1010001000000111";
			tmp(36) := "0001100000111000";
			tmp(37) := "1010001000001000";
			tmp(38) := "0001100001000011";
			tmp(39) := "1010001000001001";
			tmp(40) := "0001100000111011";
			tmp(41) := "1010001000001010";
			tmp(42) := "0001100001000001";
			tmp(43) := "1010001000001101";
			tmp(44) := "0001100001010100";
			tmp(45) := "1010001000001110";
			tmp(46) := "0001100001100111";
			tmp(47) := "1010001000001111";
			tmp(48) := "0001100001000101";
			tmp(49) := "1010001000010000";
			tmp(50) := "0001100001001000";
			tmp(51) := "1010001000010010";
			tmp(52) := "0001100001001011";
			tmp(53) := "1010001000010001";
			tmp(54) := "0001100001001110";
			tmp(55) := "0001000000001001";
			tmp(56) := "0011110000000010";
			tmp(57) := "0101101100000001";
			tmp(58) := "0001000000001001";
			tmp(59) := "0100110000000010";
			tmp(60) := "0101101100000001";
			tmp(61) := "0001000000001001";
			tmp(62) := "0100010000000010";
			tmp(63) := "0110001100000001";
			tmp(64) := "0001000000001001";
			tmp(65) := "0101010000000010";
			tmp(66) := "0001000000001001";
			tmp(67) := "0100000000001010";
			tmp(68) := "0001000000001001";
			tmp(69) := "0111110000000010";
			tmp(70) := "0111101100000001";
			tmp(71) := "0001000000001001";
			tmp(72) := "1000010000000010";
			tmp(73) := "1000001100000001";
			tmp(74) := "0001000000001001";
			tmp(75) := "1001010000000010";
			tmp(76) := "1001001100000001";
			tmp(77) := "0001000000001001";
			tmp(78) := "1000110000000000";
			tmp(79) := "1000101100000000";
		  
		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
