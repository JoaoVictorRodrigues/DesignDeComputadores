LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE dec_constants IS
    CONSTANT addr_w : NATURAL := 8;

    CONSTANT disp0 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000000";
    CONSTANT disp1 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000001";
    CONSTANT disp2 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000010";
    CONSTANT disp3 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000011";
    CONSTANT disp4 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000100";
    CONSTANT disp5 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000101";
    CONSTANT habBase : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000110";
    CONSTANT clrBase : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00000111";
    CONSTANT b3 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001000";
    CONSTANT b2 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001001";
    CONSTANT b1 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001010";
    CONSTANT b0 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001011";
    CONSTANT sw0 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001100";
    CONSTANT sw1 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001101";
    CONSTANT sw2 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001110";
    CONSTANT sw3 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00001111";
    CONSTANT sw4 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00010000";
    CONSTANT sw5 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00010001";
    CONSTANT sw6 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00010010";
    CONSTANT sw7 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00010011";
    CONSTANT sw8 : STD_LOGIC_VECTOR(addr_w - 1 DOWNTO 0) := "00010100";

END PACKAGE dec_constants;